
// 8x7 sprite memory
module letter_memory(
	input [3:0] xcoord, ycoord,
	input [3:0] letra,
	input reset,
	output Rx, Gx, Bx, on
	);
	
	localparam ROWS = 7;
	localparam WIDTH = 8;
	localparam PIXEL_WIDTH = WIDTH*3;
	
	reg [PIXEL_WIDTH-1:0] letra_mem [9:0] [ROWS-1:0];
	
	always @(posedge reset) begin
		letra_mem[0][0] <= 24'b000111111111111111000000;
		letra_mem[0][1] <= 24'b111000000000000000111000;
		letra_mem[0][2] <= 24'b111000000000000000111000;
		letra_mem[0][3] <= 24'b111000000000000000111000;
		letra_mem[0][4] <= 24'b111000000000000000111000;
		letra_mem[0][5] <= 24'b111000000000000000111000;
		letra_mem[0][6] <= 24'b000111111111111111000000;

		// Letra 1
		letra_mem[1][0] <= 24'b000111111111111000000000;
		letra_mem[1][1] <= 24'b000000000111111000000000;
		letra_mem[1][2] <= 24'b000000000111111000000000;
		letra_mem[1][3] <= 24'b000000000111111000000000;
		letra_mem[1][4] <= 24'b000000000111111000000000;
		letra_mem[1][5] <= 24'b000000000111111000000000;
		letra_mem[1][6] <= 24'b000111111111111111000000;

		// Letra 2
		letra_mem[2][0] <= 24'b000111111111111111000000;
		letra_mem[2][1] <= 24'b000000000000111111000000;
		letra_mem[2][2] <= 24'b000000000000111111000000;
		letra_mem[2][3] <= 24'b000111111111111111000000;
		letra_mem[2][4] <= 24'b000111111000000000000000;
		letra_mem[2][5] <= 24'b000111111000000000000000;
		letra_mem[2][6] <= 24'b000111111111111111000000;

		// Letra 3
		letra_mem[3][0] <= 24'b000111111111111111000000;
		letra_mem[3][1] <= 24'b000000000000111111000000;
		letra_mem[3][2] <= 24'b000000000000111111000000;
		letra_mem[3][3] <= 24'b000111111111111111000000;
		letra_mem[3][4] <= 24'b000000000000111111000000;
		letra_mem[3][5] <= 24'b000000000000111111000000;
		letra_mem[3][6] <= 24'b000111111111111111000000;
		
		// Letra 4
		letra_mem[4][0] <= 24'b000000000111111111000000;
		letra_mem[4][1] <= 24'b000000111111111111000000;
		letra_mem[4][2] <= 24'b000111111000111111000000;
		letra_mem[4][3] <= 24'b111111000000111111000000;
		letra_mem[4][4] <= 24'b111111111111111111000000;
		letra_mem[4][5] <= 24'b000000000000111111000000;
		letra_mem[4][6] <= 24'b000000000000111111000000;

		// Letra 5
		letra_mem[5][0] <= 24'b111111111111111111111000;
		letra_mem[5][1] <= 24'b111000000000000000000000;
		letra_mem[5][2] <= 24'b111000000000000000000000;
		letra_mem[5][3] <= 24'b111111111111111111111000;
		letra_mem[5][4] <= 24'b000000000000000000111000;
		letra_mem[5][5] <= 24'b000000000000000000111000;
		letra_mem[5][6] <= 24'b111111111111111111111000;

		// Letra 6
		letra_mem[6][0] <= 24'b000111111111111111000000;
		letra_mem[6][1] <= 24'b111000000000000000000000;
		letra_mem[6][2] <= 24'b111000000000000000000000;
		letra_mem[6][3] <= 24'b111111111111111111000000;
		letra_mem[6][4] <= 24'b111000000000000000111000;
		letra_mem[6][5] <= 24'b111000000000000000111000;
		letra_mem[6][6] <= 24'b000111111111111111000000;

		// Letra 7
		letra_mem[7][0] <= 24'b111111111111111111111000;
		letra_mem[7][1] <= 24'b000000000000000111111000;
		letra_mem[7][2] <= 24'b000000000000111111000000;
		letra_mem[7][3] <= 24'b000000000111111000000000;
		letra_mem[7][4] <= 24'b000000111111000000000000;
		letra_mem[7][5] <= 24'b000111111000000000000000;
		letra_mem[7][6] <= 24'b111111000000000000000000;

		// Letra 8
		letra_mem[8][0] <= 24'b000111111111111111000000;
		letra_mem[8][1] <= 24'b111000000000000000111000;
		letra_mem[8][2] <= 24'b111000000000000000111000;
		letra_mem[8][3] <= 24'b000111111111111111000000;
		letra_mem[8][4] <= 24'b111000000000000000111000;
		letra_mem[8][5] <= 24'b111000000000000000111000;
		letra_mem[8][6] <= 24'b000111111111111111000000;

		// Letra 9
		letra_mem[9][0] <= 24'b000111111111111111000000;
		letra_mem[9][1] <= 24'b111000000000000000111000;
		letra_mem[9][2] <= 24'b111000000000000000111000;
		letra_mem[9][3] <= 24'b000111111111111111111000;
		letra_mem[9][4] <= 24'b000000000000000000111000;
		letra_mem[9][5] <= 24'b000000000000000000111000;
		letra_mem[9][6] <= 24'b000111111111111111000000;	
	end

	assign Rx = letra_mem[letra][ycoord][3*(WIDTH-1-xcoord)+2];
	assign Gx = letra_mem[letra][ycoord][3*(WIDTH-1-xcoord)+1];
	assign Bx = letra_mem[letra][ycoord][3*(WIDTH-1-xcoord)+0];
	assign on = Rx == 1 && Gx == 1 && Bx == 1;

endmodule
