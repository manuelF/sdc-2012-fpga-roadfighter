
// 5x5 car sprite memory,
module car_memory(

	input [4:0] xcoord, ycoord,
	input [2:0] car,
	input reset, pclk,
//	input clk, Reset, pclk,	
	output Rx, Gx, Bx
	);
	
	
	localparam ROWS = 32;
	localparam WIDTH = 16*3;
	reg [WIDTH-1:0] carrow;
	
	reg [WIDTH-1:0] car0[ROWS-1:0]; //mi auto
	reg [WIDTH-1:0] car1[ROWS-1:0]; //auto enemigo
		
	
	// Initialize
	always @(posedge reset) 
	begin

		// Mi Auto 0
		car0[0] =  48'b111111111000000000000000000000000000000111111111;
		car0[1] =  48'b111111000000000000000000000000000000000000111111;
		car0[2] =  48'b111111000000000000000000000000000000000000111111;
		car0[3] =  48'b111111000000000000000000000000000000000000111111;
		car0[4] =  48'b111111000000000000000000000000000000000000111111;
		car0[5] =  48'b111111000000000000000000000000000000000000111111;
		car0[6] =  48'b111111000000000000000000000000000000000000111111;
		car0[7] =  48'b111111000000000000000000000000000000000000111111;
		car0[8] =  48'b111111000000000000000000000000000000000000111111;
		car0[9] =  48'b111111000000000000000000000000000000000000111111;
		car0[10] = 48'b111111000000000000000000000000000000000000111111;
		car0[11] = 48'b111111000000000000000000000000000000000000111111;
		car0[12] = 48'b111111000000000000000000000000000000000000111111;
		car0[13] = 48'b111111000000000000000000000000000000000000111111;
		car0[14] = 48'b111111000000000000000000000000000000000000111111;
		car0[15] = 48'b111111000000000000000000000000000000000000111111;
		car0[16] = 48'b111111000000000000000000000000000000000000111111;
		car0[17] = 48'b111111000000000000000000000000000000000000111111;
		car0[18] = 48'b111111000000000000000000000000000000000000111111;
		car0[19] = 48'b111111000000000000000000000000000000000000111111;
		car0[20] = 48'b111111000000000000000000000000000000000000111111;
		car0[21] = 48'b111111000000000000000000000000000000000000111111;
		car0[22] = 48'b111111000000000000000000000000000000000000111111;
		car0[23] = 48'b111111000000000000000000000000000000000000111111;
		car0[24] = 48'b111111000000000000000000000000000000000000111111;
		car0[25] = 48'b111111000000000000000000000000000000000000111111;
		car0[26] = 48'b111111000000000000000000000000000000000000111111;
		car0[27] = 48'b111111000000000000000000000000000000000000111111;
		car0[28] = 48'b111111000000000000000000000000000000000000111111;
		car0[29] = 48'b111111000000000000000000000000000000000000111111;
		car0[30] = 48'b111111000000000000000000000000000000000000111111;
		car0[31] = 48'b111111111111111111111111111111111111111111111111;

		// AutoEnemigo 1
		car1[0] =  48'b111111111000000000000000000000000000000111111111;
		car1[1] =  48'b111111000000000000000000000000000000000000111111;
		car1[2] =  48'b111111000000000000000000000000000000000000111111;
		car1[3] =  48'b111111000000000000000000000000000000000000111111;
		car1[4] =  48'b111111000000000000000000000000000000000000111111;
		car1[5] =  48'b111111000000110110110110110110110110000000111111;
		car1[6] =  48'b111111000000110110110110110110110110000000111111;
		car1[7] =  48'b111111000000110110110000000000000000000000111111;
		car1[8] =  48'b111111000000110110110000000000000000000000111111;
		car1[9] =  48'b111111000000110110110110110110110110000000111111;
		car1[10] = 48'b111111000000110110110110110110110110000000111111;
		car1[11] = 48'b111111000000110110110000000000000000000000111111;
		car1[12] = 48'b111111000000110110110000000000000000000000111111;
		car1[13] = 48'b111111000000110110110110110110110110000000111111;
		car1[14] = 48'b111111000000110110110110110110110110000000111111;
		car1[15] = 48'b111111000000000000000000000000000000000000111111;
		car1[16] = 48'b111111000000000000000000000000000000000000111111;
		car1[17] = 48'b111111000000000000000000000000000000000000111111;
		car1[18] = 48'b111111000000000000000000000000000000000000111111;
		car1[19] = 48'b111111000000000000000000000000000000000000111111;
		car1[20] = 48'b111111000000000000000000000000000000000000111111;
		car1[21] = 48'b111111000000000000000000000000000000000000111111;
		car1[22] = 48'b111111000000000000000000000000000000000000111111;
		car1[23] = 48'b111111000000000000000000000000000000000000111111;
		car1[24] = 48'b111111000000000000000000000000000000000000111111;
		car1[25] = 48'b111111000000000000000000000000000000000000111111;
		car1[26] = 48'b111111000000000000000000000000000000000000111111;
		car1[27] = 48'b111111000000000000000000000000000000000000111111;
		car1[28] = 48'b111111000000000000000000000000000000000000111111;
		car1[29] = 48'b111111000000000000000000000000000000000000111111;
		car1[30] = 48'b111111000000000000000000000000000000000000111111;
		car1[31] = 48'b111111111111111111111111111111111111111111111111;
			
	end
	/*
		return {
			ok: false
		}
		return;
		{
			ok: false;
		}
	*/
	// Assign signals to proper outputs
	/*reg R,G,B;
	always @(posedge pclk) 
	begin

		if (car == 0)
			carrow = car0[ycoord];
		if (car == 1)
			carrow = car1[ycoord];
	
		R = carrow[(xcoord*3)+2];
		G = carrow[(xcoord*3)+1];
		B = carrow[(xcoord*3)+0];		
	end
	assign Rx=R;
	assign Gx=G;
	assign Bx=B;*/
		
	
	/*
	always @(car0[0],car0[1],car0[2],car0[3],car0[4],car0[5],car0[6],car0[7],car0[8],car0[9],car0[10],car0[11],car0[12],car0[13],car0[14],car0[15],
	car0[16],car0[17],car0[18],car0[19],car0[20],car0[21],car0[22],car0[23],car0[24],car0[25],car0[26],car0[27],car0[28],car0[29],car0[30],car0[31],
car1[0],car1[1],car1[2],car1[3],car1[4],car1[5],car1[6],car1[7],car1[8],car1[9],car1[10],car1[11],car1[12],car1[13],car1[14],car1[15],
car1[16],car1[17],car1[18],car1[19],car1[20],car1[21],car1[22],car1[23],car1[24],car1[25],car1[26],car1[27],car1[28],car1[29],car1[30],car1[31]	)
	
	begin
	*/
		assign Rx = (car == 0 & car0[ycoord][(xcoord*3+2)]) | (car >= 1 & car1[ycoord][(xcoord*3)+2]);
		assign Gx = (car == 0 & car0[ycoord][(xcoord*3+1)]) | (car >= 1 & car1[ycoord][(xcoord*3)+1]);
		assign Bx = (car == 0 & car0[ycoord][(xcoord*3+0)]) | (car >= 1 & car1[ycoord][(xcoord*3)+0]);
	
/*		if(car==0)
			carrow = car0[ycoord];
		if(car>=1)
			carrow = car1[ycoord];
	//end
	assign Rx=carrow[(xcoord*3)+2];
	assign Gx=carrow[(xcoord*3)+1];
	assign Bx=carrow[(xcoord*3)+0];
	*/
endmodule